magic
tech scmos
timestamp 1710668795
<< nwell >>
rect -11 3 36 21
<< polysilicon >>
rect -5 13 -3 15
rect 0 13 2 15
rect 28 13 31 15
rect -5 2 -3 5
rect -5 -21 -3 -2
rect 0 -4 2 5
rect 28 2 31 5
rect 15 -1 31 2
rect 15 -2 18 -1
rect 4 -8 7 -5
rect 5 -21 7 -8
rect 15 -21 18 -6
rect -5 -27 -3 -25
rect 5 -27 7 -25
rect 15 -27 18 -25
<< ndiffusion >>
rect -7 -25 -5 -21
rect -3 -25 -1 -21
rect 3 -25 5 -21
rect 7 -25 9 -21
rect 13 -25 15 -21
rect 18 -25 22 -21
<< pdiffusion >>
rect -7 5 -5 13
rect -3 5 0 13
rect 2 5 7 13
rect 11 5 15 13
rect 25 5 28 13
rect 31 5 32 13
<< metal1 >>
rect -7 17 -2 21
rect 2 17 7 21
rect 11 17 25 21
rect -11 16 25 17
rect -11 13 -7 16
rect 21 13 25 16
rect -17 -2 -7 1
rect 7 0 11 5
rect 8 -3 11 0
rect -17 -8 0 -5
rect 8 -6 14 -3
rect 32 -6 36 5
rect 8 -13 11 -6
rect -1 -16 11 -13
rect 22 -10 43 -6
rect -1 -21 3 -16
rect 22 -21 26 -10
rect -11 -32 -7 -25
rect -1 -26 3 -25
rect 9 -32 13 -25
rect -11 -33 13 -32
rect -7 -37 -1 -33
rect 3 -37 9 -33
rect -11 -38 13 -37
<< ntransistor >>
rect -5 -25 -3 -21
rect 5 -25 7 -21
rect 15 -25 18 -21
<< ptransistor >>
rect -5 5 -3 13
rect 0 5 2 13
rect 28 5 31 13
<< polycontact >>
rect -7 -2 -3 2
rect 0 -8 4 -4
rect 14 -6 18 -2
<< ndcontact >>
rect -11 -25 -7 -21
rect -1 -25 3 -21
rect 9 -25 13 -21
rect 22 -25 26 -21
<< pdcontact >>
rect -11 5 -7 13
rect 7 5 11 13
rect 21 5 25 13
rect 32 5 36 13
<< psubstratepcontact >>
rect -11 -37 -7 -33
rect -1 -37 3 -33
rect 9 -37 13 -33
<< nsubstratencontact >>
rect -11 17 -7 21
rect -2 17 2 21
rect 7 17 11 21
<< labels >>
rlabel nsubstratencontact 0 19 0 19 5 Vdd
rlabel metal1 -16 -1 -16 -1 3 a
rlabel metal1 -15 -7 -15 -7 3 b
rlabel psubstratepcontact 1 -35 1 -35 1 gnd
rlabel metal1 14 -5 14 -5 7 out
rlabel metal1 39 -8 39 -8 7 ORout
<< end >>
